module nbt

#flag -I @VROOT/assets/cNBT
#include 'nbt.h'