module level

type Dimension = int

const (
	nether = Dimension(-1)
	overworld = Dimension(0)
	the_end = Dimension(1)
)