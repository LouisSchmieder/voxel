module packet

enum State {
	handshake
	status
	login
	play
}